
module Generator_reset(
input iClk,//%Input Clock
output oReset//%Output Reset
);
//////////////////////////////////////////////////////////////////////////////////
// Internal Signals
//////////////////////////////////////////////////////////////////////////////////
//!
reg [15:0] rCounter=16'h0;
reg rReset=1'b0;
//////////////////////////////////////////////////////////////////////////////////
// Continuous assignments
//////////////////////////////////////////////////////////////////////////////////
assign oReset=rReset;
//////////////////////////////////////////////////////////////////////////////////
// Sequential logic
//////////////////////////////////////////////////////////////////////////////////
always @ (posedge iClk)
	begin 
		if(rCounter != 16'h000f)
			begin		
				rCounter = rCounter+ 16'h1;
				rReset<=1'b0;
			end
		else 
			begin
				rReset<=1'b1;			
			end	 
	end
endmodule 
		
	